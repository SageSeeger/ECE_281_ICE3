library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ripple_adder_tb is
end ripple_adder_tb;

architecture test_bench of ripple_adder_tb is 
  component ripple_adder is
    Port ( A : in STD_LOGIC_VECTOR (3 downto 0);
           B : in STD_LOGIC_VECTOR (3 downto 0);
           Cin : in STD_LOGIC;
           S : out STD_LOGIC_VECTOR (3 downto 0);
           Cout : out STD_LOGIC );
  end component;
  
  signal w_addends     : std_logic_vector(7 downto 0) := x"00"; 
  signal w_sum         : std_logic_vector(3 downto 0) := x"0";
  signal w_Cin, w_Cout : std_logic;

begin
  ripple_adder_uut : ripple_adder port map (
       A    => w_addends(3 downto 0),
       B    => w_addends(7 downto 4),
       Cin  => w_Cin,
       S    => w_sum,
       Cout => w_Cout
  );
  
  test_process : process 
  begin
     -- Test all zeros input
     w_addends <= x"00"; w_Cin <= '0'; wait for 10 ns;
     assert (w_sum = x"0" and w_Cout = '0') report "bad with zeros" severity failure;

     -- Test all ones input
     w_addends <= x"FF"; w_Cin <= '1'; wait for 10 ns;
     assert (w_sum = x"F" and w_Cout = '1') report "bad with ones" severity failure;

     w_addends <= x"00"; w_Cin <= '1'; wait for 10 ns;
     assert (w_sum = x"1" and w_Cout = '0') report "bad with zero and ones" severity failure;

     w_addends <= x"45"; w_Cin <= '0'; wait for 10 ns;
     assert (w_sum = x"9" and w_Cout = '0') report "bad at 45" severity failure;

     w_addends <= x"65"; w_Cin <= '1'; wait for 10 ns;
     assert (w_sum = x"C" and w_Cout = '0') report "bad at 65 and Cin" severity failure;

     wait; -- wait forever
  end process;

end test_bench;
